// $Id: $
// File name:   sr_9bit.sv
// Created:     2/10/2016
// Author:      Vikram Manja
// Lab Section: 337-05
// Version:     1.0  Initial Design Entry
// Description: 9 bit shift register for the UART :-)
module sr_9bit
(
  input wire clk,
  input wire n_rst,
  input wire shift_strobe,
  input wire serial_in,
  output reg[7:0] packet_data,
  output reg stop_bit
);
reg[8:0] parallel_out;

flex_stp_sr 
	#(
		.NUM_BITS(9),
		.SHIFT_MSB(0)
		)
	SHIFT(
		.clk(clk),
		.n_rst(n_rst),
		.serial_in(serial_in),
		.shift_enable(shift_strobe),
		.parallel_out(parallel_out)
	);


always_comb begin
  packet_data = parallel_out[7:0];
  stop_bit = parallel_out[8];
end // end always
endmodule
