mg149@ecegrid-thin4.ecn.purdue.edu.22688:1452091460