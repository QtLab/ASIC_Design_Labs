/home/ecegrid/a/mg149/ece337/Lab2/source/tb_adder_8bit.sv