/home/ecegrid/a/mg149/ece337/Lab2/source/adder_8bit.sv